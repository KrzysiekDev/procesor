library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity control is port( 
	clk : in std_logic;
	IR : in signed(31 downto 0);
	reset : in std_logic;
	--C, Z, S,P, INT : in std_logic;
	Salu, Sbb, Sba : out signed(3 downto 0);
	Sbc : out signed(4 downto 0);
	Sid : out signed(2 downto 0);
	Sa : out signed(1 downto 0);
	Smar, Smbr, WR, RD : out std_logic
	--INTA, MIO : out bit
	);
end entity;
architecture rtl of control is 
type state_type is (fetch, fetch2, decode, MOV_R, MOV_S, ADD_R, ADD_S, SUB_R, SUB_S, LD_R, LD_S, LD_A1,LD_A2,LD_A3,LD_A4,LD_A5, CMPEQ_S, CMPEQ_A1, 
                    CMPEQ_A2, CMPEQ_A3, CMPEQ_A4, CMPEQ_A5, CMPEQ_A6, CMPGE_S, CMPGE_A1,CMPGE_A2, CMPGE_A3, CMPGE_A4, CMPGE_A5, CMPGE_A6, CMPGT_S, 
                    CMPGT_A1, CMPGT_A2, CMPGT_A3, CMPGT_A4, CMPGT_A5, CMPGT_A6, CMPLE_S, CMPLE_A1, CMPLE_A2, CMPLE_A3, CMPLE_A4, CMPLE_A5, 
                    CMPLE_A6, CMPLT_S, CMPLT_A1, CMPLT_A2, CMPLT_A3, CMPLT_A4, CMPLT_A5, CMPLT_A6, OR_S, OR_A1, OR_A2, OR_A3, OR_A4, OR_A5, OR_A6, 
                    CMPNE_R, CMPNE_S, CMPNE_A1, CMPNE_A2, CMPNE_A3, CMPNE_A4, CMPNE_A5, CMPNE_A6, BCDtoB); 
signal state : state_type;

 begin
    process (clk, reset)
        begin
            if(reset = '1') then
                state <= fetch;
            elsif (clk'event and clk = '1') then
                case state is
                    when fetch =>
                        state <= fetch2;
                    when fetch2 =>
                        state <= decode;
                    --dekodowanie rozkazu procesora
                    when decode =>
                        -- pierwsze 2 bity - ilość argumentów operacji
                        case IR(31 downto 29) is
                        	when "001" =>
                        		case IR(28 downto 26) is
                        			when "000" =>
                        				state <= BCDtoB;
                        			when others =>
                        				state <= fetch;
                        		end case;
                        	when "010" =>	
                        		case IR(28 downto 26) is
                        			when "000" => 
                        				state <= MOV_R;
                        			when "001" =>
                        				state <= ADD_R;
                        			when "010" =>
                        			 	state <= SUB_R;
                        			when "011" =>
                        			 	state <= LD_R;
                        			when "100" =>
                        			 	state <= CMPNE_R;
                        			when others =>
                        			 	state <= fetch;
                        		end case;
                        	when "011" =>
                        		case IR(28 downto 26) is
                        			when "000" => 
                        				state <= MOV_S;
                        			when "001" =>
                        				state <= ADD_S;
                        			when "010" =>
                        			 	state <= SUB_S;
                        			when others =>
                        			 	state <= fetch;
                        		end case;
                        	when "100" =>
                        		case IR(28 downto 26) is
                        			when "000" => 
                        				state <= OR_S;
                        			when others =>
                        				state <= fetch;
                        		end case;
                        	when "101" =>
                        		case IR(28 downto 26) is
                        			when "000" => 
                        				state <= LD_S;
                        			when "001" =>
                        				state <= CMPEQ_S;
                        			when "010" =>
                        			 	state <= CMPGE_S;
                        			when "011" =>
                        			 	state <= CMPGT_S;
                        			when "100" =>
                        			 	state <= CMPLE_S;
                        			when "101" =>
                        			 	state <= CMPLT_S;
                        			when "110" =>
                        			 	state <= CMPNE_S;
                        			when others =>
                        			 	state <= fetch;
                        		end case;
                        	when "110" =>
                        		case IR(28 downto 26) is
                        			when "000" => 
                        				state <= LD_A1;
                        			when "001" =>
                        				state <= CMPEQ_A1;
                        			when "010" =>
                        			 	state <= CMPGE_A1;
                        			when "011" =>
                        			 	state <= CMPGT_A1;
                        			when "100" =>
                        			 	state <= CMPLE_A1;
                        			when "101" =>
                        			 	state <= CMPLT_A1;
                        			when "110" =>
                        			 	state <= CMPNE_A1;
                                    when "111" => 
                        			     state <= OR_A1;
                                    when others =>
                        			 	state <= fetch;
                        		end case;
                        	when others =>
                        		state <= fetch;
                        end case;

                      -- przejscia pomiedzy stanami
                    when BCDtoB =>
                    	state <= fetch;
                    when MOV_R =>
                    	state <= fetch;
                    when ADD_R =>
                    	state <= fetch;
                    when SUB_R =>
                    	state <= fetch;
                    when LD_R =>
                    	state <= fetch;
                    when CMPNE_R =>
                    	state <= fetch;
                    when MOV_S =>
                    	state <= fetch;
                    when ADD_S =>
                    	state <= fetch;
                    when SUB_S =>
                    	state <= fetch;
                    when OR_S =>
                    	state <= fetch;
                    when LD_S =>
                     	state <= fetch;
                    when CMPEQ_S =>
                    	state <= fetch;
                    when CMPGE_S =>
                    	state <= fetch;
                    when CMPGT_S =>
                    	state <= fetch;
                    when CMPLE_S =>
                    	state <= fetch;
                    when CMPLT_S =>
                    	state <= fetch;
                    when CMPNE_S =>
                    	state <= fetch;
                    when LD_A1 =>
                    	state <= LD_A2;
                    when LD_A2 =>
                    	state <= LD_A3;
                    when LD_A3 =>
                    	state <= LD_A4;
                    when LD_A4 =>
                    	state <= LD_A5;
                    when LD_A5 =>
                    	state <= fetch;    
                    when CMPEQ_A1 =>
                        state <= CMPEQ_A2;
                    when CMPEQ_A2 =>
                        state <= CMPEQ_A3;
                    when CMPEQ_A3 =>
                        state <= CMPEQ_A4;
                    when CMPEQ_A4 =>
                        state <= CMPEQ_A5;
                    when CMPEQ_A5 =>
                        state <= CMPEQ_A6;
                    when CMPEQ_A6 =>
                        state <= fetch;
                    when CMPGE_A1 =>
                        state <= CMPGE_A2;
                    when CMPGE_A2 =>
                        state <= CMPGE_A3;
                    when CMPGE_A3 =>
                        state <= CMPGE_A4;
                    when CMPGE_A4 =>
                        state <= CMPGE_A5;
                    when CMPGE_A5 =>
                        state <= CMPGE_A6;
                    when CMPGE_A6 =>
                        state <= fetch;
                    when CMPGT_A1 =>
                        state <= CMPGT_A2;
                    when CMPGT_A2 =>
                        state <= CMPGT_A3;
                    when CMPGT_A3 =>
                        state <= CMPGT_A4;
                    when CMPGT_A4 =>
                        state <= CMPGT_A5;
                    when CMPGT_A5 =>
                        state <= CMPGT_A6;
                    when CMPGT_A6 =>
                        state <= fetch;
                    when CMPLE_A1 =>
                        state <= CMPLE_A2;
                    when CMPLE_A2 =>
                        state <= CMPLE_A3;
                    when CMPLE_A3 =>
                        state <= CMPLE_A4;
                    when CMPLE_A4 =>
                        state <= CMPLE_A5;
                    when CMPLE_A5 =>
                        state <= CMPLE_A6;
                    when CMPLE_A6 =>
                        state <= fetch;
                    when CMPLT_A1 =>
                        state <= CMPLT_A2;
                    when CMPLT_A2 =>
                        state <= CMPLT_A3;
                    when CMPLT_A3 =>
                        state <= CMPLT_A4;
                    when CMPLT_A4 =>
                        state <= CMPLT_A5;
                    when CMPLT_A5 =>
                        state <= CMPLT_A6;
                    when CMPLT_A6 =>
                        state <= fetch;
                    when CMPNE_A1 =>
                        state <= CMPNE_A2;
                    when CMPNE_A2 =>
                        state <= CMPNE_A3;
                    when CMPNE_A3 =>
                        state <= CMPNE_A4;
                    when CMPNE_A4 =>
                        state <= CMPNE_A5;
                    when CMPNE_A5 =>
                        state <= CMPNE_A6;
                    when CMPNE_A6 =>
                        state <= fetch;
                    when OR_A1 =>
                        state <= OR_A2;
                    when OR_A2 =>
                        state <= OR_A3;
                    when OR_A3 =>
                        state <= OR_A4;
                    when OR_A4 =>
                        state <= OR_A5;
                    when OR_A5 =>
                        state <= OR_A6;
                    when OR_A6 =>
                        state <= fetch;
                    when others =>
                    	state <= fetch;

				end case;
        	end if;
    end process;


    process(state)
    begin
    	case state is
    		when fetch =>
    			Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "01";
				Smar <= '1';
				Smbr <= '0';
				WR <= '0';
				RD <= '1';
			when fetch2 =>
				Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= "0000";
				Sid <= "001";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '1';
			when decode =>
				Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when BCDtoB =>
				Salu <="1011";
    			Sbb <= IR(3 downto 0);
    			Sbc <= "11111";
    			Sba <= IR(3 downto 0);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when MOV_R =>
				Salu <="0001";
    			Sbb <= IR(8 downto 5);
    			Sbc <= IR(4 downto 0);
    			Sba <= IR(8 downto 5);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when ADD_R =>
				Salu <="0010";
    			Sbb <= IR(8 downto 5);
    			Sbc <= IR(4 downto 0);
    			Sba <= IR(8 downto 5);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when SUB_R =>
				Salu <="0011";
    			Sbb <= IR(8 downto 5);
    			Sbc <= IR(4 downto 0);
    			Sba <= IR(8 downto 5);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when LD_R =>
				Salu <="0001";
    			Sbb <= IR(8 downto 5);
    			Sbc <= IR(4 downto 0);
    			Sba <= IR(8 downto 5);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when CMPNE_R =>
				Salu <="1010";
    			Sbb <= IR(8 downto 5);
    			Sbc <= IR(4 downto 0);
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when MOV_S =>
				Salu <="0001";
    			Sbb <= IR(15 downto 12);
    			Sbc <= "01110";
    			Sba <= IR(15 downto 12);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when ADD_S =>
				Salu <="0010";
    			Sbb <= IR(15 downto 12);
    			Sbc <= "01110";
    			Sba <= IR(15 downto 12);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when SUB_S =>
				Salu <="0011";
    			Sbb <= IR(15 downto 12);
    			Sbc <= "01110";
    			Sba <= IR(15 downto 12);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when OR_S =>
				Salu <="1001";
    			Sbb <= IR(19 downto 16);
    			Sbc <= "01111";
    			Sba <= IR(19 downto 16);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when LD_S =>
				Salu <="0001";
    			Sbb <= IR(21 downto 18);
    			Sbc <= "10000";
    			Sba <= IR(21 downto 18);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';	
			when CMPEQ_S =>
				Salu <="0100";
    			Sbb <= IR(21 downto 18);
    			Sbc <= "10000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';	
			when CMPGE_S =>
				Salu <="0101";
    			Sbb <= IR(21 downto 18);
    			Sbc <= "10000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';	
			when CMPGT_S =>
				Salu <="0110";
    			Sbb <= IR(21 downto 18);
    			Sbc <= "10000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';	
			when CMPLE_S =>
				Salu <="0111";
    			Sbb <= IR(21 downto 18);
    			Sbc <= "10000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';	
			when CMPLT_S =>
				Salu <="1000";
    			Sbb <= IR(21 downto 18);
    			Sbc <= "10000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when CMPNE_S =>
				Salu <="1010";
    			Sbb <= IR(21 downto 18);
    			Sbc <= "10000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';	
			when LD_A1 =>
				Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "01";
				Smar <= '1';
				Smbr <= '0';
				WR <= '0';
				RD <= '1';
			when LD_A2 =>
				Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= "1101";
				Sid <= "001";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when LD_A3 =>
				Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "11";
				Smar <= '1';
				Smbr <= '0';
				WR <= '0';
				RD <= '1';
			when LD_A4 =>
				Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
			when LD_A5 =>
				Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= IR(3 downto 0);
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
            when CMPEQ_A1 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "01";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPEQ_A2 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1101";
                Sid <= "001";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPEQ_A3 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "11";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPEQ_A4 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPEQ_A5 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "0001";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPEQ_A6 =>
                Salu <="0100";
                Sbb <= IR(3 downto 0);
                Sbc <= "00001";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPGE_A1 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "01";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPGE_A2 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1101";
                Sid <= "001";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPGE_A3 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "11";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPGE_A4 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPGE_A5 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "0001";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPGE_A6 =>
                Salu <="0101";
                Sbb <= IR(3 downto 0);
                Sbc <= "00001";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPGT_A1 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "01";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPGT_A2 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1101";
                Sid <= "001";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPGT_A3 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "11";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPGT_A4 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPGT_A5 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "0001";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPGT_A6 =>
                Salu <="0110";
                Sbb <= IR(3 downto 0);
                Sbc <= "00001";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPLE_A1 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "01";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPLE_A2 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1101";
                Sid <= "001";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPLE_A3 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "11";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPLE_A4 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPLE_A5 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "0001";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPLE_A6 =>
                Salu <="0111";
                Sbb <= IR(3 downto 0);
                Sbc <= "00001";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPLT_A1 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "01";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPLT_A2 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1101";
                Sid <= "001";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPLT_A3 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "11";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPLT_A4 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPLT_A5 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "0001";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPLT_A6 =>
                Salu <="1000";
                Sbb <= IR(3 downto 0);
                Sbc <= "00001";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPNE_A1 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "01";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPNE_A2 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1101";
                Sid <= "001";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPNE_A3 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "11";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when CMPNE_A4 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPNE_A5 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "0001";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when CMPNE_A6 =>
                Salu <="1010";
                Sbb <= IR(3 downto 0);
                Sbc <= "00001";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when OR_A1 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "01";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when OR_A2 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1101";
                Sid <= "001";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when OR_A3 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "11";
                Smar <= '1';
                Smbr <= '0';
                WR <= '0';
                RD <= '1';
            when OR_A4 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "1111";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when OR_A5 =>
                Salu <="0000";
                Sbb <= "0000";
                Sbc <= "00000";
                Sba <= "0001";
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
            when OR_A6 =>
                Salu <="1001";
                Sbb <= IR(3 downto 0);
                Sbc <= "00001";
                Sba <= IR(3 downto 0);
                Sid <= "000";
                Sa <= "00";
                Smar <= '0';
                Smbr <= '0';
                WR <= '0';
                RD <= '0';
			when others =>
				Salu <="0000";
    			Sbb <= "0000";
    			Sbc <= "00000";
    			Sba <= "1111";
				Sid <= "000";
				Sa <= "00";
				Smar <= '0';
				Smbr <= '0';
				WR <= '0';
				RD <= '0';
    	end case;
    end process;
end rtl;
                        	
